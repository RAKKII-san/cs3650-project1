`timescale 1 ps / 100 fs
// Verilog project: 32-bit 5-stage Pipelined MIPS Processor in Verilog 
// Shift left 2 module 
module shift_left_2(Out32, In32);
output [31:0] Out32;
input [31:0] In32;

assign Out32 = {In32[29:0],2'b00};
endmodule